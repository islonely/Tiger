module dom

// https://html.spec.whatwg.org/multipage/semantics.html#htmlheadelement
pub struct HTMLHeadElement {
	HTMLElement
}