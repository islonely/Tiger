module dom

struct EventTarget {
}