module dom

// https://html.spec.whatwg.org/multipage/grouping-content.html#htmlparagraphelement
pub struct HTMLParagraphElement {
	HTMLElement
pub mut:
	// obsolete
	align string
}