module dom

// https://html.spec.whatwg.org/multipage/grouping-content.html#htmldivelement
pub struct HTMLDivElement {
	HTMLElement
pub mut:
	// obsolete
	align string
}