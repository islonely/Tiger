module dom

// https://html.spec.whatwg.org/multipage/semantics.html#htmltitleelement
pub struct HTMLTitleElement {
	HTMLElement
pub mut:
	text string
}