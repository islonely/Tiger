module dom

pub struct Document{}