module dom

// https://html.spec.whatwg.org/multipage/media.html#htmlaudioelement
pub struct HTMLAudioElement {
	HTMLMediaElement
}
