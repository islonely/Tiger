module dom

// https://html.spec.whatwg.org/multipage/text-level-semantics.html#htmlspanelement
pub struct HTMLSpanElement {
	HTMLElement
}