module dom

// https://html.spec.whatwg.org/multipage/semantics.html#htmlhtmlelement
pub struct HTMLHtmlElement {
	HTMLElement
pub mut:
	// obsolete
	version string
}