module dom

// https://html.spec.whatwg.org/multipage/grouping-content.html#htmlmenuelement
pub struct HTMLMenuElement {
	HTMLElement
pub mut:
	// obsolete
	compact bool
}