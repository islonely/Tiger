module dom

pub struct DocumentFragment {
	Node
}