module dom

// https://html.spec.whatwg.org/multipage/edits.html#htmlmodelement
pub struct HTMLModElement {
	HTMLElement
pub mut:
	cite      string
	date_time string
}
