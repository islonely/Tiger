module components

enum VerticalAlignment {
	top
	middle
	bottom
}

enum HorizontalAlignment {
	left
	center
	right
}
