module dom

[heap]
struct Text {
	AbstractNode
}
