module dom

pub struct Element{}