module dom

// https://html.spec.whatwg.org/multipage/grouping-content.html#htmldlistelement
pub struct HTMLDListElement {
	HTMLElement
pub mut:
	compact bool
}