module dom

// https://html.spec.whatwg.org/multipage/embedded-content.html#htmlpictureelement
pub struct HTMLPictureElement {
	HTMLElement
}