module dom

// https://html.spec.whatwg.org/multipage/sections.html#htmlheadingelement
pub struct HTMLHeadingElement {
	HTMLElement
pub mut:
	// obsolete
	align string
}