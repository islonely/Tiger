module dom

pub struct HTMLAudioElement {
	HTMLMediaElement
}
