module dom

// https://html.spec.whatwg.org/multipage/grouping-content.html#htmlpreelement
pub struct HTMLPreElement {
	HTMLElement
pub mut:
	// obsolete
	width i64
}