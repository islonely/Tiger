module dom

struct EventTarget {
}
