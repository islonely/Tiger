module dom

// https://html.spec.whatwg.org/multipage/tables.html#htmltablecaptionelement
pub struct HTMLTableCaptionElement {
	HTMLElement
pub mut:
	// obsolete
	align string
}
