module dom

// https://html.spec.whatwg.org/multipage/text-level-semantics.html#htmlbrelement
pub struct HTMLBRElement {
	HTMLElement
pub mut:
	// obsolete
	clear string
}
