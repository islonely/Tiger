module dom

pub struct Comment {
	AbstractNode
__global:
	data string
}
